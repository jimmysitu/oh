module siaminer(/*AUTOARG*/);
    /*AUTOINPUT*/
    /*AUTOOUTPUT*/
    
    /*AUTOWIRE*/
    /*AUTOREG*/

    siacore uSiacore(/*AUTOINST*/);

    uart2core uUart2core(/*AUTOINST*/);
    
endmodule

