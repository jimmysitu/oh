module uartloop(/*AUTOARG*/);
    /*AUTOINPUT*/
    /*AUTOOUTPUT*/
    
    /*AUTOWIRE*/
    /*AUTOREG*/

    uart2core uUart2core(/*AUTOINST*/);
    
endmodule

